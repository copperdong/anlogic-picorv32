// Verilog netlist created by TD v3.0.987
// Thu Feb  9 11:21:40 2017

module sysmem_ml  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(14)
  (
  addra,
  cea,
  clka,
  dia,
  rsta,
  wea,
  doa
  );

  input [9:0] addra;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(19)
  input cea;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(20)
  input clka;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(21)
  input [7:0] dia;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(18)
  input rsta;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(23)
  input wea;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(22)
  output [7:0] doa;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_ml.v(16)


  AL_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0607F0260585060501F00087C78094060687F000058094470780800700000101),
    .INIT_01(256'h78E4F00087ECF00788E880FA66F08080070607F00592470F0E0E030608080505),
    .INIT_02(256'h2B722B77766A2B666650497675727266662B65706C2B656255F000F000F08760),
    .INIT_03(256'h0000000000000000000000000000000000000000003129284324462B472B2B2B),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_sub_000000_000_1024_8 (
    .addra({addra,3'b111}),
    .cea(cea),
    .clka(clka),
    .dia({open_n21,dia}),
    .rsta(rsta),
    .wea(wea),
    .doa({open_n35,doa}));

endmodule 

