// Verilog netlist created by TD v3.0.987
// Thu Feb  9 11:23:04 2017

module sysmem_hi  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(14)
  (
  addra,
  cea,
  clka,
  dia,
  rsta,
  wea,
  doa
  );

  input [9:0] addra;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(19)
  input cea;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(20)
  input clka;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(21)
  input [7:0] dia;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(18)
  input rsta;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(23)
  input wea;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(22)
  output [7:0] doa;  // /home/rgwan/anlogic/picorv32_demo/al_ip/mem_hi.v(16)


  AL_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0500FC0800110800F7FE00FFFF0000FF0000FE00000000001000001000054000),
    .INIT_01(256'hFEFEFE0000FFFC000300040302FF0000FA0510F6000200000204020204070606),
    .INIT_02(256'h2B24766674657267724832622B24676E7A756E616873714A79FC00FD01FEFFFE),
    .INIT_03(256'h00000000000000000000000000000000000000000030364E3A00514E462B2B2B),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_sub_000000_000_1024_8 (
    .addra({addra,3'b111}),
    .cea(cea),
    .clka(clka),
    .dia({open_n21,dia}),
    .rsta(rsta),
    .wea(wea),
    .doa({open_n35,doa}));

endmodule 

